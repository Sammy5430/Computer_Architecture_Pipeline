module condition_handler(output reg Cond_true, input[3:0] CC, CI, input ID_B);
	always @ (ID_B,CC,CI)
		if(ID_B)
		begin
		case(CI)
			4'b0000:
				begin
					Cond_true<=CC[2];//Z
				end
			4'b0001:
				begin
					Cond_true<=!CC[2];//~Z
				end
			4'b0010:
				begin
					Cond_true<=CC[1];//C
				end
			4'b0011:
				begin
					Cond_true<=!CC[1];//~C
				end
			4'b0100:
				begin
					Cond_true<=CC[3];//N
				end
			4'b0101:
				begin
					Cond_true<=!CC[3];//~N
				end
			4'b0110:
				begin
					Cond_true<=CC[0];//V
				end
			4'b0111:
				begin
					Cond_true<=!CC[0];//~V
				end
			4'b1000:
				begin
					Cond_true<=CC[1]&&(!CC[2]);//C&&~Z
				end
			4'b1001:
				begin
					Cond_true<=(!CC[1])||CC[2];//~C||Z
				end
			4'b1010:
				begin
					Cond_true<=CC[3]==CC[0];//N=V
				end
			4'b1011:
				begin
					Cond_true<=CC[3]!=CC[0];//N~=V
				end
			4'b1100:
				begin
					Cond_true<=(!CC[2])&&(CC[3]==CC[0]);//(~Z)&&N=V
				end
			4'b1101:
				begin
					Cond_true<=(CC[2])||(CC[3]!=CC[0]);//(Z)||N!=V
				end
			4'b1110:
				begin
					Cond_true<=1;
				end
			4'b1111:
				begin
					Cond_true<=0;
				end
		endcase
		end
		else Cond_true<=0;
endmodule		